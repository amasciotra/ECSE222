

--Alex Masciotra
--Joe Lipari

--Testbench game controller

library ieee;
library modelsim_lib;
use modelsim_lib.util.all;
use ieee.std_logic_1164.all;

-- Declare entity
entity tb_game_controller is
end tb_game_controller;

architecture behaviour of tb_game_controller is
-- Component declaration of Device Under Test (DUT)
	component game_controller is
		port (
		clk             : in std_logic; -- Clock for the system
    		rst             : in std_logic; -- Resets the state machine
    		shoot           : in std_logic; -- User shoot
		move_left       : in std_logic; -- User left
		move_right      : in std_logic; -- User right	  
		pixel_x         : in integer; -- X position of the cursor
		pixel_y		       : in integer; -- Y position of the cursor 
   	 	pixel_color	    : out std_logic_vector (2 downto 0)
   	 	
			
		);
	end component;

--Inputs
signal clk_in: std_logic;
signal rst_in: std_logic;
signal shoot_in: std_logic;
signal move_left_in : std_logic; -- User left
signal move_right_in: std_logic; -- User right		
signal move_down_in: std_logic;		  
signal pixel_x_in : integer; -- X position of the cursor
signal pixel_y_in : integer; -- Y position of the cursor  




--Outputs
signal pixel_color_out: std_logic_vector (2 downto 0);


--Helper
constant clk_period : time := 50ns;


type state is ( init, pre_game, gameplay, game_over);
signal game_state: state ;
signal lives: integer;
signal score: integer;

begin
	dut: game_controller
	port map(
		clk => clk_in,
		rst => rst_in,
		shoot => shoot_in,
		move_left =>move_left_in,
		move_right =>move_right_in,
		--move_down=>move_down_in,
		pixel_x => pixel_x_in,
		pixel_y => pixel_y_in,
		--score_temp => score_temp_in,
		--lives_temp => lives_temp_in, -- begin lives
		pixel_color => pixel_color_out
	);

	-- this process creates a clock signal
	clk_process: process
	begin
		clk_in <= '0';
		wait for clk_period/2;
		clk_in <= '1';
		wait for clk_period/2;
	end process;

	-- spy process to access signals
	spy_process: process
	begin
		init_signal_spy("/dut/current_state", "/game_state", 1);
		init_signal_spy("/dut/lives", "/lives", 1);
		init_signal_spy("/dut/score", "/score", 1);
	  wait;
	end process spy_process;

	
	-- Actual unit test
	test: process

	begin		
		pixel_x_in <= 0;
		pixel_y_in <= 0;
		shoot_in <= '0';

		rst_in <= '1';
		wait for clk_period;
		assert game_state = init report "Error: Reset does not set current state to init" severity Error;

		rst_in <= '0';
		wait for clk_period;
		assert game_state = pre_game report "Error: When init, current state does not change to pre_game" severity Error;
		
		shoot_in <= '1';
		wait for clk_period;
		assert game_state = gameplay report "Error: shooting does not start game" severity Error;
		shoot_in <= '0';
	
		--score_temp_in <= 60;
		--wait for clk_period;		
		--assert game_state = game_over report "Error: when score is 60, the game is not over" severity Error;

		shoot_in <= '1';
		wait for clk_period;
		assert game_state = init report "Error: shooting after game over does not initialize game" severity Error;
		shoot_in <= '0';
		
		assert false report "Test success!" severity failure;

	end process;

end behaviour;
